module ARM (
  input clk, rst
);


endmodule
