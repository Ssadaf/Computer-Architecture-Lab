module WB_stage (
  input clk, rst, 
  input [31:0] PC_in, 
  output [31:0] PC_out
);
  assign PC_out = PC_in;

endmodule
